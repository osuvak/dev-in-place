.tran 1.0000e-07 10m